--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Definitions is

	type EXECUTION_STATE is(	
				EXEC_STATE_READY,
				EXEC_STATE_RUNNING,
				EXEC_STATE_DONE
			 );	

end Definitions;

package body Definitions is

 
end Definitions;
