----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:03:50 02/15/2015 
-- Design Name: 
-- Module Name:    UartTransmit4Test - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity UartTransmit4Test is
	Port 
	( 
		clock : in STD_LOGIC;
		reset : in STD_LOGIC;
		RS232_dataout : out STD_LOGIC
	);
end UartTransmit4Test;

architecture Behavioral of UartTransmit4Test is

signal execution_started : std_logic;
	signal exec_done : std_logic := '0';
	signal call_1_ALU_Add_return_val : std_logic_vector(31 downto 0);
	signal call_1_ALU_Mul_return_val : std_logic_vector(31 downto 0);

	-- Serial transmission signal
	signal transmit_done : std_logic := '0';				-- Flag the entire transmission is complete
	signal transmit_started : std_logic := '0';			-- Flag to start transmission of execution data
	signal start_transmit_4bytes : std_logic := '0';	-- Flag to start transmission of 1 4byte data
	signal send_4bytes_complete : std_logic := '0';		-- Flags if the transmission of a 4byte chunk is complete
	signal data_4bytes : std_logic_vector(31 downto 0) := (others => '0'); -- 4 byte data to send 
	signal data_count : std_logic_vector(7 downto 0);

	
	component UartTransmit4 is
		Port( 
				clock : in STD_LOGIC;
				reset : in STD_LOGIC;
				start_transmit_4bytes: in STD_LOGIC;
				data_4bytes : in STD_LOGIC_VECTOR(31 downto 0);
				send_4bytes_complete : out STD_LOGIC;
				RS232_dataout : out STD_LOGIC
			 );
	end component UartTransmit4;

begin

	uart_send_4byte : UartTransmit4 port map
	(
		clock 						=> clock,
		reset 						=> reset,
		start_transmit_4bytes	=> start_transmit_4bytes,
		data_4bytes					=> data_4bytes,
		send_4bytes_complete  	=> send_4bytes_complete,
		RS232_dataout 				=> RS232_dataout
	);
	
	-- Process to transmit all data values to the serial communication device
	-- It will multiplex data values into a 4byte signal
	-- This process is generated by the compiler given all the global variable names
	proc_transmit_data : process(reset, exec_done, send_4bytes_complete)
		variable varIndex : integer := 0;
		variable canSend : boolean := false;
		
	begin
		ResetSync : if reset = '1' then
			varIndex := 0;
			canSend := false;
			data_count <= X"00";
			start_transmit_4bytes <= '0';	
			transmit_done <= '0';
			transmit_started <= '0';
			
			-- Always start for this test
			exec_done <= '1';
		
		elsif reset = '0' then
			IsExecutionDone : if exec_done = '1' then
			
				canSend := false;
				CanStartFirstTransmit : if transmit_started = '0' then
					-- Set transmit flag
					-- This controls the transmission of bits in the UartTransmit4 component
					start_transmit_4bytes <= '1'; 
					canSend := true;
				end if CanStartFirstTransmit;
				
				CanStartTransmitAfterPreviousTransmitIsDone : if send_4bytes_complete = '1' then
					canSend := true;
				end if CanStartTransmitAfterPreviousTransmitIsDone;
				
				if canSend = true then
					mux_dataval : if data_count = X"00" then
						data_4bytes <= X"41424344";
					--elsif data_count = X"01" then
					--	data_4bytes <= X"45464748";
					elsif data_count = X"01" then
						start_transmit_4bytes <= '0';
						transmit_done <= '1';
					end if mux_dataval;
				
					varIndex := to_integer(unsigned(data_count));
					varIndex := varIndex + 1;
					data_count <= std_logic_vector(to_unsigned(varIndex, 8));
					
				end if;
			end if IsExecutionDone;
		end if ResetSync;
	end process proc_transmit_data;
	

end Behavioral;

