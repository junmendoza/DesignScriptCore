
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ProgramSynthesized is
port( 
	clock : in std_logic;
	reset : in std_logic
)
end ProgramSynthesized;

architecture Behavioral of ProgramSynthesized is

signal a : std_logic_vector(31 downto 0);
signal b : std_logic_vector(31 downto 0);

begin

end Behavioral;

